

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

use work.core_pack.all;
use work.op_pack.all;

package alu_pkg is
  component alu is
    port (
  		op   : in  alu_op_type;
  		A, B : in  std_logic_vector(DATA_WIDTH-1 downto 0);
  		R    : out std_logic_vector(DATA_WIDTH-1 downto 0);
  		Z    : out std_logic;
  		V    : out std_logic
      );
  end component;
end package;


library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

use work.core_pack.all;
use work.op_pack.all;
use work.alu_pkg.all;

entity alu_tb is

end entity;

architecture alu_tb of alu_tb is

  signal op : alu_op_type;
  signal A, B : std_logic_vector(DATA_WIDTH-1 downto 0);
  signal R : std_logic_vector(DATA_WIDTH-1 downto 0);
  signal Z, V : std_logic;

begin

  test : process
  begin

  op<=alu_nop; A<="10101010010101011010101001010101"; B<="11001100001100111100110000110011"; wait for 10 ns;
  op<=alu_nop; A<="00000000000000000000000000000000"; B<="00010010001101000101011001111000"; wait for 10 ns;
  op<=alu_add; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_add; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_add; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_add; A<="00000000000000000000000000000000"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_add; A<="11111111111111111111111111111111"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_add; A<="11111111111111111111111111111111"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_add; A<="01111111111111111111111111111111"; B<="01111111111111111111111111111111"; wait for 10 ns;
  op<=alu_add; A<="10000000000000000000000000000000"; B<="10000000000000000000000000000000"; wait for 10 ns;
  op<=alu_sub; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_sub; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_sub; A<="00000000000000000000000000000000"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_sub; A<="11111111111111111111111111111111"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_sub; A<="01111111111111111111111111111111"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_sub; A<="11111111111111111111111111111110"; B<="01111111111111111111111111111111"; wait for 10 ns;
  op<=alu_and; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_and; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_or; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_or; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_or; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_xor; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_xor; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_xor; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_nor; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_nor; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_nor; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_slt; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_slt; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_slt; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_slt; A<="11111111111111111111111111111111"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_slt; A<="11111111111111111111111111111111"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_sltu; A<="00000000000000000000000000000000"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_sltu; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_sltu; A<="00000000000000000000000000000001"; B<="00000000000000000000000000000001"; wait for 10 ns;
  op<=alu_sltu; A<="00000000000000000000000000000000"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_sltu; A<="11111111111111111111111111111111"; B<="00000000000000000000000000000000"; wait for 10 ns;
  op<=alu_sltu; A<="11111111111111111111111111111111"; B<="11111111111111111111111111111111"; wait for 10 ns;
  op<=alu_sll; A<="00000000000000000000000000000100"; B<="10000111011001010100001100100001"; wait for 10 ns;
  op<=alu_sll; A<="00000000000000000000000000100100"; B<="10000111011001010100001100100001"; wait for 10 ns;
  op<=alu_srl; A<="00000000000000000000000000000100"; B<="10000111011001010100001100100001"; wait for 10 ns;
  op<=alu_srl; A<="00000000000000000000000000100100"; B<="10000111011001010100001100100001"; wait for 10 ns;
  op<=alu_sra; A<="00000000000000000000000000000100"; B<="10000111011001010100001100100001"; wait for 10 ns;
  op<=alu_sra; A<="00000000000000000000000000100100"; B<="10000111011001010100001100100001"; wait for 10 ns;
  op<=alu_lui; A<="10000111011001010100001100100001"; B<="00000000000000000000000000000000"; wait for 10 ns;



    wait;
  end process;

  alu_inst : alu
  port map (
    op => op,
    A => A,
    B => B,
    R => R,
    Z => Z,
    V => V
  );

end architecture;
