-- TODO: implement TB
